`timescale 1ns/1ps
// =============================================================================
//  Program : AGU.sv
//  Author  : Hon-Chou Dai
//  Date    : May/15/2021
// -----------------------------------------------------------------------------
//  Description:
//  Data structure used in memory opertaion.
// -----------------------------------------------------------------------------
//  Revision information:
//
//    None.
//
// -----------------------------------------------------------------------------
//  License information:
//
//  This software is released under the BSD-3-Clause Licence,
//  see https://opensource.org/licenses/BSD-3-Clause for details.
//  In the following license statements, "software" refers to the
//  "source code" of the complete hardware/software system.
//
//  Copyright 2022,
//                    Embedded Intelligent Systems Lab (EISL)
//                    Deparment of Computer Science
//                    National Yang Ming Chiao Tung Uniersity (NYCU)
//                    Hsinchu, Taiwan.
//
//  All rights reserved.
//
//  Redistribution and use in source and binary forms, with or without
//  modification, are permitted provided that the following conditions are met:
//
//  1. Redistributions of source code must retain the above copyright notice,
//     this list of conditions and the following disclaimer.
//
//  2. Redistributions in binary form must reproduce the above copyright notice,
//     this list of conditions and the following disclaimer in the documentation
//     and/or other materials provided with the distribution.
//
//  3. Neither the name of the copyright holder nor the names of its contributors
//     may be used to endorse or promote products derived from this software
//     without specific prior written permission.
//
//  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
//  AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
//  IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
//  ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
//  LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
//  CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
//  SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
//  INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
//  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
//  ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
//  POSSIBILITY OF SUCH DAMAGE.
// =============================================================================

import Falco_pkg::*;

package L1_cache_pkg;
// L1 ICache
    typedef logic [Falco_pkg::ICACHE_LINE_SIZE - 1:0] icache_line_t;
    typedef struct packed {
        Falco_pkg::mem_addr_t instr0_addr;
        Falco_pkg::mem_addr_t instr1_addr;
        logic p_strobe;
    } core_icache_req_t;

    typedef struct packed {
        Falco_pkg::raw_instruction_t raw_instr0;
        logic instr0_valid;
        Falco_pkg::raw_instruction_t raw_instr1;
        logic instr1_valid;
    } core_icache_resp_t;

    typedef struct packed {
        Falco_pkg::mem_addr_t m_addr;
        logic m_strobe;
    } icache_mem_req_t;

    typedef struct packed {
        icache_line_t m_dout;
        logic m_ready;
    } icache_mem_resp_t;

    typedef struct packed {
        logic store_req;
        Falco_pkg::mem_addr_t store_addr;
        Falco_pkg::xlen_data_t store_data;
        logic [3:0] store_mask; //byte_mask
    } core_store_req_t;

    typedef struct packed {
        logic store_finished;
        logic store_miss;
    } core_dcache_store_resp_t;

    typedef struct packed {
        logic load_req;
        Falco_pkg::mem_addr_t load_addr;
    } core_load_req_t;

    typedef struct packed {
        logic load_finished;
        logic load_miss;
        Falco_pkg::xlen_data_t load_data;
    } core_dcache_load_resp_t;
endpackage
